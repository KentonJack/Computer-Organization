module registers(clk, regwr, rreg1, rreg2, wreg, wdata, rdata1, rdata2);
	input	clk;
	input	regwr;
	input	[4:0]	rreg1, rreg2, wreg;
	input	[31:0]	wdata;
	output	[31:0]	rdata1, rdata2;
	
	reg 	[31:0]	rh[31:0];//MIPS 32??????

	initial begin			//???
/*
		rh[1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;*/
		rh[0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
/*
		rh[24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;

		rh[26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;

		rh[28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[29] = 32'b0000_0000_0000_0000_0010_1111_1111_1100;
		rh[30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		rh[31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000;*/
	end

	always @(posedge clk) begin
		if (regwr) begin
			rh[wreg] <= wdata;			//??????????
			$display(rh[10]);
		end
	end
	
	assign rdata1 = (rreg1 != 0)? rh[rreg1]:0;
	assign rdata2 = (rreg2 != 0)? rh[rreg2]:0;		//????ra?rb
endmodule
