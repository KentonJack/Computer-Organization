module datapath(clk,rst,regdst,regwr,alusrc,memwr,memtoreg,jump,branch,aluctr,rtype,extop,ins);
	input clk;
	input rst;
	input	regdst;
	input 	regwr;
	input	alusrc;
	input	memwr;
	input	memtoreg;
	input	jump;
	input 	extop;
	input	branch;
	input [2:0]	aluctr;
	input 	rtype;
	wire [31:0] pc_now;
	wire [31:0] pc_temp;
	wire [31:0] pc_next;
	wire [31:0] pc_4;
	wire [31:0] pc_br;			//pc??,??pc???????
	wire [4:0] wreg;			//??????????
	wire [31:0] rdata1;
	wire [31:0] rdata2;
	wire [31:0] const_or_addr;
	wire [31:0] busa;
	wire [31:0] busb;
	wire zero;
	wire [31:0] aluresult;
	wire [31:0] rdata;
	wire [31:0] wdata;
	output [31:0] ins;		//???????
	pc pcgo(clk,rst,pc_next,pc_now);	//pc
	assign pc_4 = pc_now + 4;
	alu pc_alu(.busa(pc_4),.busb({const_or_addr[29:0],2'b00}),.aluctr(3'b000),.result(pc_br));
	mux2 #(32) br_mux(pc_4,pc_br,(branch & zero),pc_temp);			//???pc_4??pc_br
	mux2 #(32) j_mux(pc_temp,{pc_4[31:28],ins[25:0],2'b00},jump,pc_next);	//????????????,?????pc_next???????????
	im_4k im(pc_now[11:2],ins);		//??pc???????
	mux2 #(5) wreg_mux(ins[20:16],ins[15:11],regdst,wreg);			//??regdst???????????????rd??rt
	registers register(clk,regwr,ins[25:21],ins[20:16],wreg,wdata,rdata1,rdata2);
	ext ext(ins[15:0],extop,const_or_addr);			//????????
	assign busa = rdata1;					//busa??
	mux2 #(32) alusrc_mun(rdata2,const_or_addr,alusrc,busb);		//busb??
	//aluctrl aluctrl2(aluop,ins[5:0],rtype,aluctr);		//alu??????alu?????
	alu alu2(busa,busb,aluctr,zero,aluresult);		//alu??
	dm_4k dm(.addr(aluresult),.datain(rdata2),.memwr(memwr),.clk(clk),.dout(rdata));	//????????(alu??????????????????,busB????????,????????,clk,?????)
	mux2 #(32) regsrc_mux(aluresult,rdata,memtoreg,wdata);		//???alu???????????????wdata????????
endmodule
