 module cpu(clk,rst);
	input clk;
	input rst;
	wire [31:0] ins;		//??
	wire regdst;			//R?????????
	wire regwr;			//R?????????????????
	wire memwr;			//??????????
	wire alusrc;			//???busB???????alu??????
	wire memtoreg;			//?????alu?????????????????????
	wire jump;			//???????
	wire branch;			//???????
	wire rtype;			//???r???
	wire extop;			//????????
	wire [2:0] aluctr;		//
	control control(ins[31:26],regdst,regwr,alusrc,memwr,memtoreg,jump,branch,aluctr,rtype,extop);		//??????
	datapath datapath(clk,rst,regdst,regwr,alusrc,memwr,memtoreg,jump,branch,aluctr,rtype,extop,ins);	//???????????????????????????????????
endmodule

